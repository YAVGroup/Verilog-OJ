module top_module(
  output out
);
  // Write your code here
endmodule